`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name:full_sub
//////////////////////////////////////////////////////////////////////////////////


module full_sub (D, Bin, Bout, A, B);
    input A, B, Bin; 
	output Bout, D;

	assign D = A ^ B ^ Bin;
	assign Bout = (~A & (B^Bin)) | (B & Bin);
         
endmodule