`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name: out_reg
// By Kushalta Paudel
//////////////////////////////////////////////////////////////////////////////////

module out_reg (
    input clk_in, rst, outR, outCarry
    
	output reg 
    );   



	
	always @(posedge clk_in)
		if(rst)
			begin
				
				
			end
		else
			begin
				
			end	

endmodule  